module types

pub type PathImageOnServer = string
