module interfaces

pub interface IProfileService {
	contain(uuid string) bool
}
