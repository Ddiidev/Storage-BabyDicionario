module ws

import veb

pub struct Context {
	veb.Context
}
