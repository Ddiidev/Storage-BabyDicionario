module types

pub type PathAudioOnServer = string
